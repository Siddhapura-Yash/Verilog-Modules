// AND Gate Implementation
module and_gate(a, b, y);

input a, b;  // Inputs
output y;    // Output

assign y = a & b;  // AND operation

endmodule
