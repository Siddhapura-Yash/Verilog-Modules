// XOR Gate Implementation
module xor_gate(a, b, y);

input a, b;  // Inputs
output y;    // Output

assign y = a ^ b;  // XOR operation

endmodule
