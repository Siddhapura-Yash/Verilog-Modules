// NOT Gate Implementation
module not_gate(a, y);

input a;  // Input
output y; // Output

assign y = ~a;  // NOT operation

endmodule
